magic
tech sky130A
timestamp 1634664404
<< nwell >>
rect -45 135 200 275
<< nmos >>
rect -80 0 -65 100
rect 115 0 130 100
<< pmos >>
rect 75 155 90 255
rect 115 155 130 255
<< ndiff >>
rect -130 85 -80 100
rect -130 15 -120 85
rect -95 15 -80 85
rect -130 0 -80 15
rect -65 85 -15 100
rect -65 15 -55 85
rect -30 15 -15 85
rect -65 0 -15 15
rect 65 85 115 100
rect 65 15 75 85
rect 100 15 115 85
rect 65 0 115 15
rect 130 85 180 100
rect 130 15 140 85
rect 165 15 180 85
rect 130 0 180 15
<< pdiff >>
rect 25 240 75 255
rect 25 170 40 240
rect 65 170 75 240
rect 25 155 75 170
rect 90 155 115 255
rect 130 240 180 255
rect 130 170 140 240
rect 165 170 180 240
rect 130 155 180 170
<< ndiffc >>
rect -120 15 -95 85
rect -55 15 -30 85
rect 75 15 100 85
rect 140 15 165 85
<< pdiffc >>
rect 40 170 65 240
rect 140 170 165 240
<< psubdiff >>
rect -180 85 -130 100
rect -180 15 -165 85
rect -140 15 -130 85
rect -180 0 -130 15
rect 15 85 65 100
rect 15 15 30 85
rect 55 15 65 85
rect 15 0 65 15
<< nsubdiff >>
rect -25 240 25 255
rect -25 170 -10 240
rect 15 170 25 240
rect -25 155 25 170
<< psubdiffcont >>
rect -165 15 -140 85
rect 30 15 55 85
<< nsubdiffcont >>
rect -10 170 15 240
<< poly >>
rect 220 315 260 325
rect 220 310 230 315
rect 75 295 230 310
rect 250 295 260 315
rect 75 255 90 295
rect 220 285 260 295
rect 115 255 130 270
rect 75 130 90 155
rect -80 115 90 130
rect 115 130 130 155
rect 220 135 260 145
rect 220 130 230 135
rect 115 115 230 130
rect 250 115 260 135
rect -80 100 -65 115
rect 115 100 130 115
rect 220 105 260 115
rect -80 -15 -65 0
rect 115 -15 130 0
<< polycont >>
rect 230 295 250 315
rect 230 115 250 135
<< locali >>
rect 220 315 310 325
rect 220 295 230 315
rect 250 305 310 315
rect 250 295 260 305
rect 220 285 260 295
rect -20 245 70 250
rect -20 170 -10 245
rect 15 170 40 245
rect 65 170 70 245
rect -20 160 70 170
rect 135 240 175 250
rect 135 170 140 240
rect 165 170 175 240
rect 135 160 175 170
rect 220 135 310 145
rect 220 115 230 135
rect 250 125 310 135
rect 250 115 260 125
rect 220 105 260 115
rect -175 85 -85 95
rect -175 15 -165 85
rect -140 15 -120 85
rect -95 15 -85 85
rect -175 5 -85 15
rect -60 85 -20 95
rect -60 15 -55 85
rect -30 15 -20 85
rect -60 5 -20 15
rect 20 85 110 95
rect 20 15 30 85
rect 55 15 75 85
rect 100 15 110 85
rect 20 5 110 15
rect 135 85 175 95
rect 135 15 140 85
rect 165 15 175 85
rect 135 5 175 15
<< viali >>
rect -10 240 15 245
rect -10 175 15 240
rect 40 240 65 245
rect 40 175 65 240
rect 140 170 165 240
rect -165 15 -140 85
rect -120 15 -95 85
rect -55 15 -30 85
rect 30 15 55 85
rect 75 15 100 85
rect 140 15 165 85
<< metal1 >>
rect -15 255 70 305
rect -20 245 70 255
rect -20 175 -10 245
rect 15 175 40 245
rect 65 175 70 245
rect -20 165 70 175
rect 135 240 175 250
rect 135 170 140 240
rect 165 170 175 240
rect 135 150 175 170
rect -180 130 175 150
rect -180 125 -20 130
rect -175 85 -85 95
rect -175 15 -165 85
rect -140 15 -120 85
rect -95 15 -85 85
rect -175 5 -85 15
rect -60 85 -20 125
rect -60 15 -55 85
rect -30 15 -20 85
rect -60 5 -20 15
rect 20 85 110 95
rect 20 15 30 85
rect 55 15 75 85
rect 100 15 110 85
rect 20 5 110 15
rect 135 85 175 130
rect 135 15 140 85
rect 165 15 175 85
rect 135 5 175 15
rect -105 -30 -85 5
rect 90 -30 110 5
rect -105 -45 110 -30
<< labels >>
rlabel metal1 -180 135 -180 135 7 VOUT
port 1 e
rlabel locali 310 315 310 315 3 A
port 2 w
rlabel locali 310 135 310 135 3 B
port 3 w
rlabel metal1 25 305 25 305 1 VDD
port 4 n
rlabel metal1 -10 -45 -10 -45 5 GND
port 5 s
<< end >>
