magic
tech sky130A
timestamp 1634626743
<< nwell >>
rect -120 135 85 275
<< nmos >>
rect 0 0 15 100
<< pmos >>
rect 0 155 15 255
<< ndiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 85 65 100
rect 15 15 30 85
rect 50 15 65 85
rect 15 0 65 15
<< pdiff >>
rect -50 240 0 255
rect -50 170 -35 240
rect -15 170 0 240
rect -50 155 0 170
rect 15 240 65 255
rect 15 170 30 240
rect 50 170 65 240
rect 15 155 65 170
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
<< pdiffc >>
rect -35 170 -15 240
rect 30 170 50 240
<< psubdiff >>
rect -100 85 -50 100
rect -100 15 -85 85
rect -60 15 -50 85
rect -100 0 -50 15
<< nsubdiff >>
rect -100 240 -50 255
rect -100 170 -85 240
rect -60 170 -50 240
rect -100 155 -50 170
<< psubdiffcont >>
rect -85 15 -60 85
<< nsubdiffcont >>
rect -85 170 -60 240
<< poly >>
rect 0 255 15 270
rect 0 100 15 155
rect 0 -15 15 0
rect -25 -25 15 -15
rect -25 -45 -15 -25
rect 5 -45 15 -25
rect -25 -55 15 -45
<< polycont >>
rect -15 -45 5 -25
<< locali >>
rect -95 240 -5 250
rect -95 170 -85 240
rect -60 170 -35 240
rect -15 170 -5 240
rect -95 160 -5 170
rect 20 240 60 250
rect 20 170 30 240
rect 50 170 60 240
rect 20 160 60 170
rect 40 95 60 160
rect -95 85 -5 95
rect -95 15 -85 85
rect -60 15 -35 85
rect -15 15 -5 85
rect -95 5 -5 15
rect 20 85 60 95
rect 20 15 30 85
rect 50 15 60 85
rect 20 5 60 15
rect 40 -15 60 5
rect -100 -25 15 -15
rect -100 -35 -15 -25
rect -25 -45 -15 -35
rect 5 -45 15 -25
rect 40 -35 90 -15
rect -25 -55 15 -45
<< viali >>
rect -85 170 -60 240
rect -35 170 -15 240
rect -85 15 -60 85
rect -35 15 -15 85
<< metal1 >>
rect -120 240 85 250
rect -120 170 -85 240
rect -60 170 -35 240
rect -15 170 85 240
rect -120 160 85 170
rect -120 85 85 95
rect -120 15 -85 85
rect -60 15 -35 85
rect -15 15 85 85
rect -120 5 85 15
<< end >>
